// --------------------------------------------------------------------
// Copyright (c) 2011 by Terasic Technologies Inc. 
// --------------------------------------------------------------------
//
//
// --------------------------------------------------------------------
//
// Major Functions:	G Sensor utilization
//
// --------------------------------------------------------------------
//
// Revision History :
// --------------------------------------------------------------------
//   Ver  :| Author              :| Mod. Date   :| Changes Made:
//   V1.0 :| Rosaline Lin        :| 02/16/2011  :| Initial Revision
// --------------------------------------------------------------------

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module GSensorPose(
    iClk50Mhz,
	 iRst_n,
	 
	 iDataX,
	 iDataXVal,

	 oPosDval,
	 oXpos
 
);

//=======================================================
//  PARAMETER declarations
//=======================================================
`include "spi_param.h"

//=======================================================
//  PORT declarations
//=======================================================

input 			iClk50Mhz;
input 			iRst_n;
	 
input	[15:0]	iDataX;
input        	iDataXVal;

output reg	      oPosDval;
output reg [31:0] oXpos;

//=======================================================
//  REG/WIRE declarations
//=======================================================
 reg signed [31:0]  rVelX, rVelY, rVelZ;
 reg signed [31:0]  rPosX, rPosY, rPosZ;
 reg signed [31:0]  rDeltaVelX, rDeltaVelY, rDeltaVelZ;
 reg signed [15:0]  rAccX, rAccY, rAccZ;
 reg [31:0]  rTimeX, rTimeY, rTimeZ;
 reg signed [31:0]  rTimeCounter, rTimeCounter_d;
 reg [2:0]   rPoseState;
//=======================================================
//  Structural coding
//=======================================================
 wire 	wClk1us;
Clkdiv #( .CLKFREQ(50000000), .EXCEPTCLK(1_000_000), .multipleX(4) ) U_Clk1us
        (   
            .iClk50M(iClk50Mhz), // 50Mhz clock 
            .iRst_n(iRst_n),
//            .oError(oLEDG[0]),  // if CLKFREQ/2 great than ExpectClk, you will get a error
//            .oSampClk(oSampClk),  // multipleX expect clock, for SignalTap use
            .oClk(wClk1us)     // ExpectClk clock
        );
 
 reg rPreDataXVal1us, rPreClk1us;
  always@(posedge iClk50Mhz or negedge iRst_n) begin
     if(!iRst_n) begin
	      rTimeCounter <= 0;  rPreDataXVal1us <= 0; rPreClk1us <= 0;
	  end else begin
	  	   rPreDataXVal1us <= iDataXVal;
			rPreClk1us <= wClk1us;
			
			if( {rPreDataXVal1us, iDataXVal} == 2'b01 ) begin
				 rTimeCounter <= 0;
			end else if({rPreClk1us, wClk1us} ==2'b01)begin
			    rTimeCounter <= rTimeCounter +1;
			end
			else begin
			    rTimeCounter <= rTimeCounter;
			end
	  end
 end
 
 reg     rPreDataXVal;
 always@(posedge iClk50Mhz or negedge iRst_n) begin
     if(!iRst_n) begin
	      rVelX <= 0; rVelY <= 0; rVelZ <=0;
			rAccX <= 0; rAccY <= 0; rAccZ <= 0;
	      rTimeX <= 0; rTimeY <= 0; rTimeZ <=0;
			rPreDataXVal <= 0;  rPoseState <= 0; rTimeCounter_d <= 0;
	  end else begin
	  	   rVelX <= rVelX; rVelY <= rVelY; rVelZ <=rVelZ; 
			rAccX <= rAccX;
	      rTimeX <= rTimeX; rTimeY <= rTimeX; rTimeZ <=rTimeX;
			rPreDataXVal <= rPreDataXVal; rPoseState <= rPoseState;
			oPosDval <= 0; oXpos <= oXpos;
			/* ========================== */
         rTimeCounter_d <= rTimeCounter;
			case (rPoseState)
				0: begin
					rPreDataXVal <= iDataXVal;
					if( {rPreDataXVal, iDataXVal}==2'b01 ) begin
						rTimeX <= rTimeCounter_d;
						rAccX <= iDataX;
						rPoseState <= 1;
					end 
				end
				1: begin
				  rVelX <= rVelX + rAccX * 980* rTimeX; /* unit cm/s */
				  rPoseState <= 2;
				end
				2: begin
				  oXpos <= oXpos + rVelX * rTimeX; /* x coordinator unit cm */
				  oPosDval <= 1;
				  rPoseState <= 0;
				end
			
			endcase
			
	  end
 end

endmodule

