// --------------------------------------------------------------------
// Copyright (c) 2011 by Terasic Technologies Inc. 
// --------------------------------------------------------------------
//
// Permission:
//
// --------------------------------------------------------------------
//
// Major Functions:	G Sensor utilization
//
// --------------------------------------------------------------------
//
// Revision History :
// --------------------------------------------------------------------
//   Ver  :| Author              :| Mod. Date   :| Changes Made:
//   V1.0 :| Rosaline Lin        :| 02/16/2011  :| Initial Revision
// --------------------------------------------------------------------

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE0_NANO_G_Sensor(

    //////////// CLOCK //////////
    CLOCK_50,

    //////////// LED //////////
    LED,

    //////////// KEY //////////
    KEY,

    //////////// Accelerometer and EEPROM //////////
    G_SENSOR_CS_N,
    G_SENSOR_INT,
    I2C_SCLK,
    I2C_SDAT,
    GPIO
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input                       CLOCK_50;

//////////// LED //////////
output           [7:0]      LED;

//////////// KEY //////////
input            [1:0]      KEY;

//////////// Accelerometer and EEPROM //////////
output                      G_SENSOR_CS_N;
input                       G_SENSOR_INT;
output                      I2C_SCLK;
inout                       I2C_SDAT;
output  [35:0]              GPIO;
//=======================================================
//  REG/WIRE declarations
//=======================================================
wire                        dly_rst;
wire                        spi_clk, spi_clk_out;
wire    [15:0]              data_x;
wire                        wRst_n;
//=======================================================
//  Structural coding
//=======================================================
assign wRst_n = KEY[0];

DataCalcRate u_DataCalcRate(
                 .iClk50M(CLOCK_50),
                 .iRst_n(wRst_n),
                 
                 .iDataValid(wDvalX),
                 .oDataRateSec(GPIO),
                 
                 );

//  重置模塊
//  這個模塊負責產生一個延遲的重置信號
reset_delay u_reset_delay( 
            .iRSTN(wRst_n),          // 從按鍵0接收重置信號
            .iCLK(CLOCK_50),         // 50MHz的時鐘輸入
            .oRST(dly_rst));         // 輸出延遲的重置信號


//  初始設置和數據讀回模塊
//  這個模塊負責配置SPI並讀回數據
wire   [15:0]  wDataX, wDataY, wDataZ;
wire           wDvalX;
spi_ee_config u_spi_ee_config (
                        .iClk50M        (CLOCK_50),
                        .iRst_n          (!dly_rst),             // 使用反向的延遲重置信號
                        .iG_INT2        (G_SENSOR_INT),         // G感測器的中斷信號輸入
                        .oAcc_X         (wDataX),
                        .oAcc_Y         (wDataY),
                        .oAcc_Z         (wDataZ),
                        .oAccDval       (wDvalX),
                        /* SPI 3-wires */
                        .SPI_SDIO       (I2C_SDAT),            // SPI的雙向數據線
                        .oSPI_CSN       (G_SENSOR_CS_N),       // SPI的片選信號輸出
                        .oSPI_CLK       (I2C_SCLK));           // SPI的時鐘輸出

// LED驅動模塊
// 這個模塊負責驅動LED顯示
led_driver u_led_driver	( 
                        .iRSTN  (!dly_rst),             // 使用反向的延遲重置信號
                        .iCLK   (CLOCK_50),             // 50MHz的時鐘輸入
                        .iDIG   (wDataX[9:0]),          // 10位的數據輸入
                        .iG_INT2(wDvalX),               // G感測器的中斷信號輸入
                        .oLED   (LED));                 // LED輸出


GSensorPose GSensorPose(
    .iClk50Mhz (CLOCK_50),
     .iRst_n    (!dly_rst),
     
     .iDataX    (wDataX),
     .iDataXVal (wDvalX),

     .oPosDval  (),
     .oXpos     ()
 
);
endmodule
